package alu_pkg;
  `include "trans.sv"
  `include "gen.sv"
  `include "drv.sv"
  `include "mon.sv"
  `include "ref.sv"
  `include "sb.sv"
  `include "env.sv"
  `include "test.sv"
endpackage
