`timescale 1ns/1ns
`define op_len     8
`define cmd_len     4
`define no_of_transactions 50
